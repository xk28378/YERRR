-- Created by @(#)$CDS: vhdlin version 6.1.7-64b 09/27/2016 19:46 (sjfhw304) $
-- on Thu Oct 21 17:13:06 2021


architecture structural of inverter is

begin
      output7 <= not input7;
end structural;
