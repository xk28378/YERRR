-- Created by @(#)$CDS: vhdlin version 6.1.7-64b 09/27/2016 19:46 (sjfhw304) $
-- on Thu Oct 21 17:12:32 2021


architecture structural of and2 is

begin

  output <= input1 and input2;

end structural;
