-- Created by @(#)$CDS: vhdlin version 6.1.7-64b 09/27/2016 19:46 (sjfhw304) $
-- on Mon Nov 29 23:10:23 2021


library STD;
library IEEE;                      
use IEEE.std_logic_1164.all;       

entity tran_gate is                      
  port ( sel   : in std_logic;
         input : in std_logic;
         output:out std_logic);
end tran_gate;                          
