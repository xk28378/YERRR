-- Created by @(#)$CDS: vhdlin version 6.1.7-64b 09/27/2016 19:46 (sjfhw304) $
-- on Thu Oct 21 17:13:06 2021


library STD;
library IEEE;
use IEEE.std_logic_1164.all;

entity inverter is
	port (
		input7 : in std_logic;
		output7: out std_logic);
end inverter;
