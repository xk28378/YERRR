-- Created by @(#)$CDS: vhdlin version 6.1.7-64b 09/27/2016 19:46 (sjfhw304) $
-- on Thu Nov 18 11:10:58 2021


library STD;
library IEEE;
use IEEE.std_logic_1164.all;

entity mux_2_1 is port (
  in1: in std_logic;
  in2: in std_logic;
  sel: in std_logic;
  out1: out std_logic);
end mux_2_1;
